//parameter declaration
//FIFO
parameter X2P_SFIFO_AW_DATA_WIDTH = 56;
parameter X2P_SFIFO_AR_DATA_WIDTH = 56;
parameter X2P_SFIFO_WD_DATA_WIDTH = 36;
parameter X2P_SFIFO_RD_DATA_WIDTH = 42;
parameter POINTER_WIDTH           = 4;

//parameter SLAVE_NUM is used to set number of APB slave

//address of Register block
parameter A_START_REG     = 32'h0000_0000;
parameter A_END_REG       = 32'h0000_0FFF; 
//address of SLAVE APB
parameter A_START_SLAVE0  = 32'h0000_1000;
parameter A_END_SLAVE0    = 32'h0000_1FFF;
parameter A_START_SLAVE1  = 32'h0000_2000;
parameter A_END_SLAVE1    = 32'h0000_2FFF;
parameter A_START_SLAVE2  = 32'h0000_3000;
parameter A_END_SLAVE2    = 32'h0000_3FFF;
parameter A_START_SLAVE3  = 32'h0000_4000;
parameter A_END_SLAVE3    = 32'h0000_4FFF;
parameter A_START_SLAVE4  = 32'h0000_5000;
parameter A_END_SLAVE4    = 32'h0000_5FFF;
parameter A_START_SLAVE5  = 32'h0000_6000;
parameter A_END_SLAVE5    = 32'h0000_6FFF;
parameter A_START_SLAVE6  = 32'h0000_7000;
parameter A_END_SLAVE6    = 32'h0000_7FFF;
parameter A_START_SLAVE7  = 32'h0000_8000;
parameter A_END_SLAVE7    = 32'h0000_8FFF;
parameter A_START_SLAVE8  = 32'h0000_9000;
parameter A_END_SLAVE8    = 32'h0000_9FFF;
parameter A_START_SLAVE9  = 32'h0000_A000;
parameter A_END_SLAVE9    = 32'h0000_AFFF;
parameter A_START_SLAVE10 = 32'h0000_B000;
parameter A_END_SLAVE10   = 32'h0000_BFFF;
parameter A_START_SLAVE11 = 32'h0000_C000;
parameter A_END_SLAVE11   = 32'h0000_CFFF;
parameter A_START_SLAVE12 = 32'h0000_D000;
parameter A_END_SLAVE12   = 32'h0000_DFFF;
parameter A_START_SLAVE13 = 32'h0000_E000;
parameter A_END_SLAVE13   = 32'h0000_EFFF;
parameter A_START_SLAVE14 = 32'h0000_F000;
parameter A_END_SLAVE14   = 32'h0000_FFFF;
parameter A_START_SLAVE15 = 32'h0001_0000;
parameter A_END_SLAVE15   = 32'h0001_0FFF;
parameter A_START_SLAVE16 = 32'h0001_1000;
parameter A_END_SLAVE16   = 32'h0001_1FFF;
parameter A_START_SLAVE17 = 32'h0001_2000;
parameter A_END_SLAVE17   = 32'h0001_2FFF;
parameter A_START_SLAVE18 = 32'h0000_3000;
parameter A_END_SLAVE18   = 32'h0001_3FFF;
parameter A_START_SLAVE19 = 32'h0001_4000;
parameter A_END_SLAVE19   = 32'h0001_4FFF;
parameter A_START_SLAVE20 = 32'h0001_5000;
parameter A_END_SLAVE20   = 32'h0001_5FFF;
parameter A_START_SLAVE21 = 32'h0001_6000;
parameter A_END_SLAVE21   = 32'h0001_6FFF;
parameter A_START_SLAVE22 = 32'h0001_7000;
parameter A_END_SLAVE22   = 32'h0001_7FFF;
parameter A_START_SLAVE23 = 32'h0001_8000;
parameter A_END_SLAVE23   = 32'h0001_8FFF;
parameter A_START_SLAVE24 = 32'h0001_9000;
parameter A_END_SLAVE24   = 32'h0001_9FFF;
parameter A_START_SLAVE25 = 32'h0001_A000;
parameter A_END_SLAVE25   = 32'h0001_AFFF;
parameter A_START_SLAVE26 = 32'h0001_B000;
parameter A_END_SLAVE26   = 32'h0001_BFFF;
parameter A_START_SLAVE27 = 32'h0001_C000;
parameter A_END_SLAVE27   = 32'h0001_CFFF;
parameter A_START_SLAVE28 = 32'h0001_D000;
parameter A_END_SLAVE28   = 32'h0001_DFFF;
parameter A_START_SLAVE29 = 32'h0001_E000;
parameter A_END_SLAVE29   = 32'h0001_EFFF;
parameter A_START_SLAVE30 = 32'h0001_F000;
parameter A_END_SLAVE30   = 32'h0001_FFFF;
parameter A_START_SLAVE31 = 32'h0002_0000;
parameter A_END_SLAVE31   = 32'h0002_0FFF;